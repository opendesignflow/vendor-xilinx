module b ;


endmodule
