`include "defs.h"
`include "test.h"
module a ;
    
    reg t [`SIZE:0];
     
    b b_I();

endmodule
